module state_timer (
        input rst_n,    // Active low asynchronous clock
        input clk,      // System clock
);
        
endmodule